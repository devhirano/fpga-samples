module whitespace2(
    a,
    b,
    c,
    y,
    z);

input a;
input b;
input c;
output y;
output z;

wire a;
wire b;
wire c;
wire y;
wire z;

endmodule
