// this is comment
/* this is comment */

module hello;

initial begin
    $display ("Hello World");
    #10 $finish;
end

endmodule
