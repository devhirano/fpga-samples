module comment(a,b,c,y,z);

/*
multi
line
comment
*/

// single line comment

input a,b,c;  // comment after impl
output y,z;

wire a,b,c;
reg y,z;


endmodule
