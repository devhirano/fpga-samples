module whitespace1(a,b,c,y,z);
input a,b,c; output y,z;
wire a,b,c,y,z; endmodule
