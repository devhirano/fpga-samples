module main;
  initial 
    begin
      $display("Hello, Wolrd");
      $finish;
    end
endmodule
