module numbers;

reg[31:0] one;

initial begin
    one = 1
    $display ("one = %h", one);
end

endmodule

